	--  ############ Insert Only the Usefor Sections ################


---------- DEFAULT LIBRARY ---------
library IEEE;
	use IEEE.STD_LOGIC_1164.all;
	use IEEE.NUMERIC_STD.ALL;
--	use IEEE.MATH_REAL.all;
------------------------------------
	
	
---------- OTHERS LIBRARY ----------
-- NONE
------------------------------------




entity GenricVHDL is
	generic(

		--------- SECTION ----------
		-- NONE
		----------------------------

	);
	port ( 

		--------- SECTION ----------
		-- NONE
		----------------------------	

	);                                 
end GenricVHDL;

architecture Behavioral of GenricVHDL is


	------------------ CONSTANT DECLARATION -------------------------
	
	--------- SECTION ----------
	-- NONE
	----------------------------
	
	-----------------------------------------------------------------

	
	
	------------------------ TYPES DECLARATION ----------------------

	--------- SECTION ----------
	-- NONE
	----------------------------	
	
	-----------------------------------------------------------------		

	
	
	--------------------- FUNCTIONS DECLARATION ---------------------

	--------- SECTION ----------
	-- NONE
	----------------------------	
	
	-----------------------------------------------------------------		

	
	
	
	--------------------- COMPONENTS DECLARETION --------------------

	----- First Component-------
	----------------------------	

	
	----- Last Component--------
	----------------------------	
	
	-----------------------------------------------------------------
	



	---------------------------- SIGNALS ----------------------------

	------- First Signals-------
	-- NONE
	----------------------------	

	------- Last Signals--------
	-- NONE
	----------------------------	

	--------- SECTION ----------
	-- NONE
	----------------------------
	
	----------------------------------------------------------------




	-------------------------- ATTRIBUTES --------------------------

	--------- SECTION ----------
	-- NONE
	----------------------------	
	
	-----------------------------------------------------------------

	


begin


	--------------------- COMPONENTS INSTANTIATIONS -------------------
	
	----- First Component-------
	-- NONE
	----------------------------	

	
	----- Last Component--------
	-- NONE
	----------------------------	

	
	-------------------------------------------------------------------


	
	----------------------------- DATA FLOW ---------------------------
	
	--------- SECTION ----------
	-- NONE
	----------------------------
	
	-------------------------------------------------------------------



	----------------------------- PROCESS ------------------------------

	------ Sync Process --------
	-- NONE
	----------------------------	

	
	----- Async Process --------
	-- NONE
	----------------------------


	--------- SECTION ----------
	-- NONE
	----------------------------	
	
	-------------------------------------------------------------------


end Behavioral;

